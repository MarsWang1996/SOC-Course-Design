library verilog;
use verilog.vl_types.all;
entity tb_Sobel_enhancement is
end tb_Sobel_enhancement;
